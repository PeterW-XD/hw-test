`timescale 1ns/100ps
module audio_tb;

logic clk;
logic read;
logic write;
logic [2:0] address;
logic SD;
logic SCK;
logic WS;
logic reset;
logic [31:0]readdata, writedata;
logic irq;
//logic [13:0] fft_real, fft_imag;

audio audio_init(	
	.clk(clk),	// 50M, 20ns
	.reset(reset),
	.chipselect(1'd1),
	.read(read),
	.write(write),
	.writedata(writedata),
	.address(address),
	.SD1(SD),
	.SD2(),
	.SD3(),
	.SCK(SCK),	// Sampling rate * 32 bits * 2 channels: 325ns
	
	.WS(WS),		// Smapling rate * 2 channels,
	.irq(irq),
	.readdata(readdata)
	);

always #10 clk = ~clk;
always #160 SCK = ~SCK;

// 4157 lines		
initial begin
clk = 0;
SCK = 0;
SD = 0;
address = 0;
read = 0;
write = 0;
writedata = 0;
reset = 1;
@(posedge clk) reset = 0;


//
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(posedge clk) write = 1; address = 0; writedata = 0;
@(posedge clk)	address = 1; writedata = 1;
@(posedge clk) write = 1; address = 0; writedata = 0;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk)	write = 0; address = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

#62000
@(posedge clk) write = 1; read = 0; address = 0; writedata = 0;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 1;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 2;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 3;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 4;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 5;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 6;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 7;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 8;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 9;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 10;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 11;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 12;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 13;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 14;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 15;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 16;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 17;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 18;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 19;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 20;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 21;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 22;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 23;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 24;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 25;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 26;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 27;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 28;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 29;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 30;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 31;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 32;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 33;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 34;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 35;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 36;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 37;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 38;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 39;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 40;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 41;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 42;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 43;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 44;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 45;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 46;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 47;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 48;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 49;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 50;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 51;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 52;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 53;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 54;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 55;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 56;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 57;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 58;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 59;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 60;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 61;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 62;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 63;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 64;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 65;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 66;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 67;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 68;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 69;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 70;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 71;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 72;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 73;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 74;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 75;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 76;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 77;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 78;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 79;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 80;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 81;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 82;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 83;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 84;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 85;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 86;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 87;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 88;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 89;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 90;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 91;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 92;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 93;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 94;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 95;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 96;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 97;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 98;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 99;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 100;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 101;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 102;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 103;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 104;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 105;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 106;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 107;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 108;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 109;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 110;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 111;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 112;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 113;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 114;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 115;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 116;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 117;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 118;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 119;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 120;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 121;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 122;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 123;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 124;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 125;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 126;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 127;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 128;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 129;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 130;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 131;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 132;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 133;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 134;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 135;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 136;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 137;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 138;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 139;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 140;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 141;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 142;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 143;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 144;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 145;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 146;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 147;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 148;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 149;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 150;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 151;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 152;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 153;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 154;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 155;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 156;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 157;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 158;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 159;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 160;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 161;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 162;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 163;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 164;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 165;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 166;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 167;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 168;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 169;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 170;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 171;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 172;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 173;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 174;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 175;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 176;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 177;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 178;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 179;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 180;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 181;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 182;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 183;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 184;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 185;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 186;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 187;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 188;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 189;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 190;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 191;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 192;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 193;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 194;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 195;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 196;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 197;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 198;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 199;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 200;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 201;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 202;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 203;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 204;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 205;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 206;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 207;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 208;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 209;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 210;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 211;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 212;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 213;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 214;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 215;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 216;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 217;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 218;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 219;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 220;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 221;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 222;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 223;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 224;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 225;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 226;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 227;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 228;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 229;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 230;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 231;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 232;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 233;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 234;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 235;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 236;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 237;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 238;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 239;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 240;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 241;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 242;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 243;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 244;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 245;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 246;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 247;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 248;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 249;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 250;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 251;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 252;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 253;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 254;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 255;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 256;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 257;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 258;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 259;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 260;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 261;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 262;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 263;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 264;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 265;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 266;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 267;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 268;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 269;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 270;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 271;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 272;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 273;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 274;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 275;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 276;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 277;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 278;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 279;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 280;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 281;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 282;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 283;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 284;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 285;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 286;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 287;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 288;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 289;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 290;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 291;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 292;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 293;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 294;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 295;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 296;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 297;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 298;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 299;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 300;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 301;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 302;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 303;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 304;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 305;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 306;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 307;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 308;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 309;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 310;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 311;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 312;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 313;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 314;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 315;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 316;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 317;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 318;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 319;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 320;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 321;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 322;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 323;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 324;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 325;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 326;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 327;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 328;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 329;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 330;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 331;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 332;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 333;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 334;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 335;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 336;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 337;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 338;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 339;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 340;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 341;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 342;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 343;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 344;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 345;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 346;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 347;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 348;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 349;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 350;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 351;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 352;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 353;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 354;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 355;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 356;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 357;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 358;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 359;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 360;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 361;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 362;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 363;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 364;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 365;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 366;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 367;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 368;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 369;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 370;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 371;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 372;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 373;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 374;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 375;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 376;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 377;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 378;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 379;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 380;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 381;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 382;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 383;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 384;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 385;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 386;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 387;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 388;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 389;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 390;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 391;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 392;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 393;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 394;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 395;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 396;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 397;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 398;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 399;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 400;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 401;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 402;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 403;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 404;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 405;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 406;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 407;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 408;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 409;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 410;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 411;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 412;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 413;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 414;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 415;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 416;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 417;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 418;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 419;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 420;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 421;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 422;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 423;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 424;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 425;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 426;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 427;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 428;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 429;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 430;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 431;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 432;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 433;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 434;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 435;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 436;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 437;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 438;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 439;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 440;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 441;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 442;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 443;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 444;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 445;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 446;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 447;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 448;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 449;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 450;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 451;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 452;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 453;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 454;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 455;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 456;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 457;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 458;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 459;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 460;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 461;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 462;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 463;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 464;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 465;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 466;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 467;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 468;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 469;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 470;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 471;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 472;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 473;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 474;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 475;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 476;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 477;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 478;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 479;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 480;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 481;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 482;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 483;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 484;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 485;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 486;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 487;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 488;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 489;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 490;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 491;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 492;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 493;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 494;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 495;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 496;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 497;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 498;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 499;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 500;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 501;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 502;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 503;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 504;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 505;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 506;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 507;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 508;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 509;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 510;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 511;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 512;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 513;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 514;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 515;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 516;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 517;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 518;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 519;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 520;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 521;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 522;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 523;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 524;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 525;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 526;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 527;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 528;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 529;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 530;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 531;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 532;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 533;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 534;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 535;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 536;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 537;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 538;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 539;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 540;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 541;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 542;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 543;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 544;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 545;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 546;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 547;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 548;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 549;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 550;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 551;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 552;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 553;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 554;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 555;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 556;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 557;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 558;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 559;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 560;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 561;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 562;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 563;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 564;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 565;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 566;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 567;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 568;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 569;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 570;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 571;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 572;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 573;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 574;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 575;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 576;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 577;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 578;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 579;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 580;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 581;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 582;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 583;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 584;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 585;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 586;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 587;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 588;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 589;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 590;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 591;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 592;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 593;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 594;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 595;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 596;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 597;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 598;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 599;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 600;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 601;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 602;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 603;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 604;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 605;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 606;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 607;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 608;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 609;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 610;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 611;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 612;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 613;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 614;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 615;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 616;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 617;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 618;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 619;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 620;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 621;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 622;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 623;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 624;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 625;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 626;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 627;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 628;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 629;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 630;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 631;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 632;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 633;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 634;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 635;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 636;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 637;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 638;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 639;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 640;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 641;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 642;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 643;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 644;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 645;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 646;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 647;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 648;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 649;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 650;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 651;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 652;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 653;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 654;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 655;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 656;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 657;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 658;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 659;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 660;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 661;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 662;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 663;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 664;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 665;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 666;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 667;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 668;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 669;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 670;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 671;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 672;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 673;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 674;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 675;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 676;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 677;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 678;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 679;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 680;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 681;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 682;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 683;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 684;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 685;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 686;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 687;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 688;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 689;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 690;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 691;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 692;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 693;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 694;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 695;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 696;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 697;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 698;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 699;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 700;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 701;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 702;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 703;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 704;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 705;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 706;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 707;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 708;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 709;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 710;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 711;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 712;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 713;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 714;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 715;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 716;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 717;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 718;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 719;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 720;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 721;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 722;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 723;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 724;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 725;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 726;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 727;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 728;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 729;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 730;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 731;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 732;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 733;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 734;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 735;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 736;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 737;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 738;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 739;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 740;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 741;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 742;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 743;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 744;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 745;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 746;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 747;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 748;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 749;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 750;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 751;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 752;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 753;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 754;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 755;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 756;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 757;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 758;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 759;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 760;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 761;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 762;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 763;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 764;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 765;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 766;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 767;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 768;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 769;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 770;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 771;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 772;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 773;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 774;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 775;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 776;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 777;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 778;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 779;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 780;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 781;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 782;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 783;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 784;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 785;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 786;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 787;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 788;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 789;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 790;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 791;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 792;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 793;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 794;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 795;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 796;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 797;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 798;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 799;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 800;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 801;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 802;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 803;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 804;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 805;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 806;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 807;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 808;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 809;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 810;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 811;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 812;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 813;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 814;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 815;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 816;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 817;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 818;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 819;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 820;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 821;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 822;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 823;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 824;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 825;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 826;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 827;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 828;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 829;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 830;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 831;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 832;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 833;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 834;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 835;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 836;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 837;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 838;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 839;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 840;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 841;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 842;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 843;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 844;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 845;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 846;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 847;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 848;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 849;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 850;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 851;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 852;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 853;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 854;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 855;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 856;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 857;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 858;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 859;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 860;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 861;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 862;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 863;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 864;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 865;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 866;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 867;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 868;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 869;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 870;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 871;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 872;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 873;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 874;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 875;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 876;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 877;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 878;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 879;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 880;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 881;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 882;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 883;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 884;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 885;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 886;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 887;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 888;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 889;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 890;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 891;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 892;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 893;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 894;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 895;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 896;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 897;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 898;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 899;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 900;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 901;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 902;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 903;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 904;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 905;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 906;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 907;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 908;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 909;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 910;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 911;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 912;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 913;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 914;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 915;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 916;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 917;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 918;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 919;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 920;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 921;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 922;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 923;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 924;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 925;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 926;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 927;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 928;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 929;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 930;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 931;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 932;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 933;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 934;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 935;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 936;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 937;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 938;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 939;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 940;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 941;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 942;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 943;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 944;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 945;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 946;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 947;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 948;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 949;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 950;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 951;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 952;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 953;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 954;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 955;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 956;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 957;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 958;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 959;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 960;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 961;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 962;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 963;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 964;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 965;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 966;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 967;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 968;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 969;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 970;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 971;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 972;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 973;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 974;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 975;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 976;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 977;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 978;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 979;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 980;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 981;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 982;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 983;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 984;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 985;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 986;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 987;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 988;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 989;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 990;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 991;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 992;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 993;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 994;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 995;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 996;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 997;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 998;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 999;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 1000;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 1001;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 1002;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 1003;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 1004;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 1005;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 1006;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 1007;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 1008;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 1009;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 1010;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 1011;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 1012;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 1013;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 1014;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 1015;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 1016;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 1017;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 1018;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 1019;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 1020;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 1021;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 1022;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;
@(posedge clk) write = 1; read = 0; address = 0; writedata = 1023;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk) write = 0; read = 1; address = 0;

@(posedge clk) read = 0; address = 0;

$stop;
end

endmodule