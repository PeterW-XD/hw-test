`timescale 1ns/100ps
module audio_tb;

logic clk;
logic read;
logic write;
logic [2:0] address;
logic SD;
logic SCK;
logic WS;
logic reset;
logic [31:0]readdata, writedata;
logic irq;
//logic [13:0] fft_real, fft_imag;

audio audio_init(	
	.clk(clk),	// 50M, 20ns
	.reset(reset),
	.chipselect(1'd1),
	.read(read),
	.write(write),
	.writedata(writedata),
	.address(address),
	.SD1(SD),
	.SD2(),
	.SD3(),
	.SCK(SCK),	// Sampling rate * 32 bits * 2 channels: 325ns
	
	.WS(WS),		// Smapling rate * 2 channels,
	.irq(irq),
	.readdata(readdata)
	);

always #10 clk = ~clk;
always #160 SCK = ~SCK;

// 4157 lines		
initial begin
clk = 0;
SCK = 0;
SD = 0;
address = 0;
read = 0;
write = 0;
writedata = 0;
reset = 1;
@(posedge clk) reset = 0;


//
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(posedge clk) write = 1; address = 0; writedata = 0;
@(posedge clk)	address = 1; writedata = 1;
@(posedge clk) write = 1; address = 0; writedata = 0;
@(posedge clk) address = 1; writedata = 0;
@(posedge clk)	write = 0; address = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)

@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK) SD = 0;
@(negedge SCK) SD = 1;
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)
@(negedge SCK)



#70000


$stop;
end

endmodule